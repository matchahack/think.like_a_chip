module glitchable_password_led (
    input  wire        clk,
    input  wire [7:0]  password_input,
    input  wire        button_1,   // "Enter"
    input  wire        button_0,   // Glitch or reset
    output logic [2:0] led
);

// === Parameters === //
localparam [7:0] SECRET_PASSWORD = 8'b11000111;  // 0xC7
localparam integer BLINK_PERIOD = 6_000_000;    // ~0.5 sec at 48 MHz (adjust as needed)
localparam integer DELAY_PER_BIT = 16'd1024;

// === FSM === //
typedef enum logic [1:0] {
    IDLE,
    CHECKING,
    SUCCESS,
    FAIL
} state_t;

state_t state = IDLE;

// === Registers === //
logic [2:0]  check_index;
logic [15:0] bit_delay_counter;
logic [31:0] counter;
logic reset_sync;
logic [24:0] blink_counter;
logic blink_on;

// === Reset sync === //
always_ff @(posedge clk) begin
    reset_sync <= (state == IDLE && button_0);
end

// === Main FSM === //
always_ff @(posedge clk) begin
    if (reset_sync) begin
        state             <= IDLE;
        check_index       <= 0;
        counter           <= 0;
        bit_delay_counter <= 0;
        blink_counter     <= 0;
        blink_on          <= 0;
        led               <= 3'b111;
    end else begin
        case (state)
            IDLE: begin
                led               <= 3'b111;
                counter           <= 0;
                check_index       <= 0;
                bit_delay_counter <= 0;
                blink_counter     <= 0;
                blink_on          <= 0;
                if (button_1) state <= CHECKING;
            end

            CHECKING: begin
                // Blink visible RED during checking period
                if (blink_counter < BLINK_PERIOD) begin
                    blink_counter <= blink_counter + 1;
                    blink_on      <= 1;
                    led           <= 3'b110; // RED
                end else begin
                    blink_counter <= 0;
                    blink_on      <= 0;
                    led           <= 3'b000;

                    // After visible blink, do the actual comparison
                    if (check_index < 8) begin
                        if (password_input[check_index] == SECRET_PASSWORD[check_index]) begin
                            check_index <= check_index + (button_0 ? 2 : 1);  // glitchable jump
                        end else begin
                            state <= FAIL;
                        end
                    end else begin
                        state <= SUCCESS;
                    end
                end
            end

            SUCCESS: begin
                counter <= counter + 1;
                case (counter)
                    0           : led <= 3'b110; // RED
                    30_000_000  : led <= 3'b011; // BLUE
                    60_000_000  : led <= 3'b101; // GREEN
                    default: begin end
                endcase
            end

            FAIL: begin
                led <= 3'b000;
                if (!button_1) state <= IDLE;
            end
        endcase
    end
end

endmodule
